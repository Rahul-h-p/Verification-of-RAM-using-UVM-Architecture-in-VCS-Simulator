
	class ram_virtual_sequencer extends uvm_sequencer #(uvm_sequence_item) ;
   
	`uvm_component_utils(ram_virtual_sequencer)

	ram_wr_sequencer wr_seqrh[];
	ram_rd_sequencer rd_seqrh[];
	

  	ram_env_config m_cfg;


 	extern function new(string name = "ram_virtual_sequencer",uvm_component parent);
	extern function void build_phase(uvm_phase phase);
	endclass

	function ram_virtual_sequencer::new(string name="ram_virtual_sequencer",uvm_component parent);
		super.new(name,parent);
	endfunction

	function void ram_virtual_sequencer::build_phase(uvm_phase phase);
	  if(!uvm_config_db #(ram_env_config)::get(this,"","ram_env_config",m_cfg))
		`uvm_fatal("CONFIG","cannot get() m_cfg from uvm_config_db. Have you set() it?")
    		 super.build_phase(phase);

wr_seqrh=new[m_cfg.no_of_duts];
rd_seqrh=new[m_cfg.no_of_duts];
    		
	endfunction
