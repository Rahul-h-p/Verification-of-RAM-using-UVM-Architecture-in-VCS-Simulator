

class ram_env_config extends uvm_object;


bit has_functional_coverage = 0;
bit has_wagent_functional_coverage = 0;
bit has_scoreboard = 1;
bit has_wagent = 1;
bit has_ragent = 1;
bit has_virtual_sequencer = 1;

ram_wr_agent_config m_wr_agent_cfg[];
ram_rd_agent_config m_rd_agent_cfg[];

int no_of_duts;

`uvm_object_utils(ram_env_config)

extern function new(string name = "ram_env_config");

endclass: ram_env_config

function ram_env_config::new(string name = "ram_env_config");
  super.new(name);
endfunction


