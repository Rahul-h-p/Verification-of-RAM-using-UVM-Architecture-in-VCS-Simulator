
	class ram_rd_agt_top extends uvm_env;

	`uvm_component_utils(ram_rd_agt_top)
    
      	 ram_rd_agent agnth;

	extern function new(string name = "ram_rd_agt_top" , uvm_component parent);
	extern function void build_phase(uvm_phase phase);
	extern task run_phase(uvm_phase phase);
  endclass

   	function ram_rd_agt_top::new(string name = "ram_rd_agt_top" , uvm_component parent);
		super.new(name,parent);
	endfunction

    
       	function void ram_rd_agt_top::build_phase(uvm_phase phase);
     		super.build_phase(phase);
   		agnth=ram_rd_agent::type_id::create("agnth",this);
	endfunction


	task ram_rd_agt_top::run_phase(uvm_phase phase);
		uvm_top.print_topology;
	endtask   


